module systolic_array (
    north_0_in, north_1_in, north_2_in, north_3_in,
    west_0_in, west_1_in, west_2_in, west_3_in,
);
    
endmodule